module sample();

endmodule
